// Pre-defined MACROS
`define DEPTH 8
`define WIDTH 16

